// Decodificador com base no livro de Idoeta
module DecodificadorDecimalDisplay7Seg(
    input  [3:0] I,           // 4 bits de entrada
    output a, b, c, d, e, f, g // segmentos do display
);

    // Faz wires no input
    wire A, B, C, D;

    // Faz tipo um destructuring, melhor que usar I[0], I[1]
    assign {A, B, C, D} = I;

    // -------------------------
    // Segmento a - acende para: 0,2,3,5,6,7,8,9
    // -------------------------
    assign a = ~(
          (~A & ~B & ~C & ~D) |  // 0000 - 0
          (~A & ~B &  C & ~D) |  // 0010 - 2
          (~A & ~B &  C &  D) |  // 0011 - 3
          (~A &  B & ~C &  D) |  // 0101 - 5
          (~A &  B &  C & ~D) |  // 0110 - 6
          (~A &  B &  C &  D) |  // 0111 - 7
          ( A & ~B & ~C & ~D) |  // 1000 - 8
          ( A & ~B & ~C &  D)    // 1001 - 9
    );

    // -------------------------
    // Segmento b - acende para: 0,1,2,3,4,7,8,9
    // -------------------------
    assign b = ~(
          (~A & ~B & ~C & ~D) |  // 0000 - 0
          (~A & ~B & ~C &  D) |  // 0001 - 1
          (~A & ~B &  C & ~D) |  // 0010 - 2
          (~A & ~B &  C &  D) |  // 0011 - 3
          (~A &  B & ~C & ~D) |  // 0100 - 4
          (~A &  B &  C &  D) |  // 0111 - 7
          ( A & ~B & ~C & ~D) |  // 1000 - 8
          ( A & ~B & ~C &  D)    // 1001 - 9
    );

    // -------------------------
    // Segmento c - acende para: 0,1,3,4,5,6,7,8,9
    // -------------------------
    assign c = ~(
          (~A & ~B & ~C & ~D) |  // 0000 - 0
          (~A & ~B & ~C &  D) |  // 0001 - 1
          (~A & ~B &  C &  D) |  // 0011 - 3
          (~A &  B & ~C & ~D) |  // 0100 - 4
          (~A &  B & ~C &  D) |  // 0101 - 5
          (~A &  B &  C & ~D) |  // 0110 - 6
          (~A &  B &  C &  D) |  // 0111 - 7
          ( A & ~B & ~C & ~D) |  // 1000 - 8
          ( A & ~B & ~C &  D)    // 1001 - 9
    );

    // -------------------------
    // Segmento d - acende para: 0,2,3,5,6,8,9
    // -------------------------
    assign d = ~(
          (~A & ~B & ~C & ~D) |  // 0000 - 0
          (~A & ~B &  C & ~D) |  // 0010 - 2
          (~A & ~B &  C &  D) |  // 0011 - 3
          (~A &  B & ~C &  D) |  // 0101 - 5
          (~A &  B &  C & ~D) |  // 0110 - 6
          ( A & ~B & ~C & ~D) |  // 1000 - 8
          ( A & ~B & ~C &  D)    // 1001 - 9
    );

    // -------------------------
    // Segmento e - acende para: 0,2,6,8
    // -------------------------
    assign e = ~(
          (~A & ~B & ~C & ~D) |  // 0000 - 0
          (~A & ~B &  C & ~D) |  // 0010 - 2
          (~A &  B &  C & ~D) |  // 0110 - 6
          ( A & ~B & ~C & ~D)    // 1000 - 8
    );

    // -------------------------
    // Segmento f - acende para: 0,4,5,6,8,9
    // -------------------------
    assign f = ~(
          (~A & ~B & ~C & ~D) |  // 0000 - 0
          (~A &  B & ~C & ~D) |  // 0100 - 4
          (~A &  B & ~C &  D) |  // 0101 - 5
          (~A &  B &  C & ~D) |  // 0110 - 6
          ( A & ~B & ~C & ~D) |  // 1000 - 8
          ( A & ~B & ~C &  D)    // 1001 - 9
    );

    // -------------------------
    // Segmento g - acende para: 2,3,4,5,6,8,9
    // -------------------------
    assign g = ~(
          (~A & ~B &  C & ~D) |  // 0010 - 2
          (~A & ~B &  C &  D) |  // 0011 - 3
          (~A &  B & ~C & ~D) |  // 0100 - 4
          (~A &  B & ~C &  D) |  // 0101 - 5
          (~A &  B &  C & ~D) |  // 0110 - 6
          ( A & ~B & ~C & ~D) |  // 1000 - 8
          ( A & ~B & ~C &  D)    // 1001 - 9
    );

endmodule
